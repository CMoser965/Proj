/*
Author: Christian Moser
Date: 10-28-2022
Project Description:

Create floating-point multiplier used for MLP neural network implementation.
*/

module multiplier(clk, rst, x, w, carry);

