module tanh #(N = 32)
(
    input   [N-1:0] in;
    output  [N-1:0] out;
);

endmodule